// RUN: python3 $LAKEROAD_DIR/bin/convert_module_to_btor.py \
// RUN:   --top counter --infile %s 2>/dev/null \
// RUN:   | FileCheck %s

module counter(input clk, input rst, output [7:0] out);
  logic [7:0] counter_reg;
  logic [7:0] counter_incremented;

  assign counter_incremented = counter_reg + 8'b1;
  assign out = counter_reg;

  initial begin
    counter_reg = 8'b0;
  end

  always @ (posedge clk) begin
    if (rst) counter_reg <= 8'b0;
    else counter_reg <= counter_incremented;
  end
endmodule

// CHECK: ; BTOR description generated by Yosys
// CHECK: 1 sort bitvec 1
// CHECK: 2 input 1 clk
// CHECK: 3 input 1 rst
// CHECK: 4 sort bitvec 8
// CHECK: 5 const 4 00000000
// CHECK: 6 state 4
// CHECK: 7 init 4 6 5
// CHECK: 8 state 4
// CHECK: 9 init 4 8 5
// CHECK: 10 const 1 1
// CHECK: 11 state 1
// CHECK: 12 init 1 11 10
// CHECK: 13 sort bitvec 2
// CHECK: 14 concat 13 2 11
// CHECK: 15 const 13 10
// CHECK: 16 eq 1 14 15
// CHECK: 17 ite 4 16 8 6
// CHECK: 18 output 17 out
// CHECK: 19 uext 4 10 7
// CHECK: 20 add 4 17 19
// CHECK: 21 uext 4 20 0 counter_incremented
// CHECK: 22 uext 4 17 0 counter_reg
// CHECK: 23 next 4 6 17
// CHECK: 24 ite 4 3 5 20
// CHECK: 25 next 4 8 24
// CHECK: 26 next 1 11 2
// CHECK: ; end of yosys output