module impl(input [15:0] a, b, output [15:0] o);
  assign o = a * b;
endmodule